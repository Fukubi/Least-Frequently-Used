library verilog;
use verilog.vl_types.all;
entity tb_lfu is
end tb_lfu;
